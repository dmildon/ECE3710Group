module tb_RegFile_Alu ();

endmodule
