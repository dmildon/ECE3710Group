module RegFile ();

endmodule 


