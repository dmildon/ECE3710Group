module CPU ();

endmodule
