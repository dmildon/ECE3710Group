module Register ();

endmodule
