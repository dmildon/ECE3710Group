module ALU ()

endmodule 

